module top(DA, AA, BA, MB, FS, SS, SA, MD, RW, CONSTANT, DATA);







endmodule
