module RegisterFile(index, val);
	input [2:0] index;
	output [15:0] val;







endmodule
