module RegisterFile (index, val);
	input [2:0] index;
	output [7:0] val;

	reg [7:0] register [0:15];








endmodule
